module BancoDeRegistradores();
	
	
endmodule