module Processador(b);
	output b;
	assign b = 1;
	
endmodule