module ULA();

endmodule